--------------------------------------------------------------------------------
-- Author:        {user.name} ({user.email})
--
-- Create Date:   {time:"%d-%m-%Y"}
-- Module Name:   {file}
--------------------------------------------------------------------------------
